module Two_to_one_MUX_tb; 
reg [31:0] A, B;
reg sel;
wire [31:0] out;

Two_to_one_MUX myMUX(.sel(sel), .A(A), .B(B), .out(out));

initial begin
  A = 32'b00000000000000000000000000000000;
  B = 32'b00000000000000000000000000000000;
  sel = 0;
  #100 B = 32'b00000000000000000000000000000001;
  #100 A = 32'b00000000000000000000000000000010; B = 32'b00000000000000000000000000000100;
  #100 B = 32'b00000000000000000000000000000001;
  
  #100 A = 32'b00000000000000000000000000010000; B = 32'b00000000000000000000000000000000;
  #100 sel = 1; 
  #100 B = 32'b00000000000000000000000000000001;
  #100 A = 32'b00000000000000000000000000000010; B = 32'b00000000000000000000000000000100;
  #100 B = 32'b00000000000000000000000000001000;

  
   #100 $finish;  //stop simulation
end

initial
  $monitor(
    "sel=%b A=%b B=%b out=%b",
    sel, A, B, out);

endmodule
