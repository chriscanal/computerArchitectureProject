module regFile (readAddress0, readAddress1, writeAddress, writeData, writeEnable, clk, readData0, readData1);
  input [4:0] readAddress0, readAddress1, writeAddress;
  input [31:0] writeData;
  input writeEnable, clk;
  output reg [31:0] readData0, readData1;

  reg [31:0] rF [31:0];

  initial //Set register to hold all 0s
  begin
    rF[5'b00000] = 32'b00000000000000000000000000000000;
    rF[5'b00001] = 32'b00000000000000000000000000000000;
    rF[5'b00010] = 32'b00000000000000000000000000000000;
    rF[5'b00011] = 32'b00000000000000000000000000000000;
    rF[5'b00100] = 32'b00000000000000000000000000000000;
    rF[5'b00101] = 32'b00000000000000000000000000000000;
    rF[5'b00110] = 32'b00000000000000000000000000000000;
    rF[5'b00111] = 32'b00000000000000000000000000000000;
    rF[5'b01000] = 32'b00000000000000000000000000000000;
    rF[5'b01001] = 32'b00000000000000000000000000000000;
    rF[5'b01010] = 32'b00000000000000000000000000000000;
    rF[5'b01011] = 32'b00000000000000000000000000000000;
    rF[5'b01100] = 32'b00000000000000000000000000000000;
    rF[5'b01101] = 32'b00000000000000000000000000000000;
    rF[5'b01110] = 32'b00000000000000000000000000000000;
    rF[5'b01111] = 32'b00000000000000000000000000000000;
    rF[5'b10000] = 32'b00000000000000000000000000000000;
    rF[5'b10001] = 32'b00000000000000000000000000000000;
    rF[5'b10010] = 32'b00000000000000000000000000000000;
    rF[5'b10011] = 32'b00000000000000000000000000000000;
    rF[5'b10100] = 32'b00000000000000000000000000000000;
    rF[5'b10101] = 32'b00000000000000000000000000000000;
    rF[5'b10110] = 32'b00000000000000000000000000000000;
    rF[5'b10111] = 32'b00000000000000000000000000000000;
    rF[5'b11000] = 32'b00000000000000000000000000000000;
    rF[5'b11001] = 32'b00000000000000000000000000000000;
    rF[5'b11010] = 32'b00000000000000000000000000000000;
    rF[5'b11011] = 32'b00000000000000000000000000000000;
    rF[5'b11100] = 32'b00000000000000000000000000000000;
    rF[5'b11101] = 32'b00000000000000000000000000000000;
    rF[5'b11110] = 32'b00000000000000000000000000000000;
    rF[5'b11111] = 32'b00000000000000000000000000000000;
  end
  
  always @ (readAddress0 or readAddress1)
    begin
      readData0 = rF[readAddress0];
      readData1 = rF[readAddress1];
    end

  always @ (posedge clk)
    begin
      if (writeEnable)
	rF[writeAddress] = writeData;
    end

endmodule


